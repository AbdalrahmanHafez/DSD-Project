library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity acc is
	port (
		clk				: IN STD_LOGIC;
		GSENSOR_CS_N	: OUT STD_LOGIC;
		GSENSOR_INT1	: IN STD_LOGIC;
		GSENSOR_INT2 	: IN STD_LOGIC;
		GSENSOR_SCLK 	: OUT STD_LOGIC;
		GSENSOR_SDI 	: BUFFER STD_LOGIC_VECTOR(15 downto 0);
		GSENSOR_SDO 	: BUFFER STD_LOGIC;
		sevenseg1		: OUT STD_LOGIC_VECTOR(7 downto 0);
		sevenseg2		: OUT STD_LOGIC_VECTOR(7 downto 0)
	);
end entity acc;


architecture arc_acc of acc is
	
begin
	GSENSOR_CS_N <= '0';
	GSENSOR_SDO <= '0';
	GSENSOR_SCLK<= clk;
	sevenseg1 <= "10011110";
	
	process
	begin
		wait until clk'EVENT and clk ='1';
		sevenseg2 <= "11001100";

	end process;

end architecture arc_acc;